library verilog;
use verilog.vl_types.all;
entity tb_ALU is
end tb_ALU;
